library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity REGISTRO_ESTADO is
    Port ( banderas_in : in  STD_LOGIC_VECTOR (3 downto 0);
           LF : in  STD_LOGIC;
           clr : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           banderas_out : out  STD_LOGIC_VECTOR (3 downto 0));
end REGISTRO_ESTADO;

architecture REGISTRO_ESTADO_ARCH of REGISTRO_ESTADO is

begin

	process(clk, clr)
	begin
		if(clr = '1') then
			banderas_out <= (others => '0');
		elsif(falling_edge(clk)) then
			if(LF = '1') then
				banderas_out <= banderas_in;
			end if;
		end if;
	end process;

end REGISTRO_ESTADO_ARCH;

